library verilog;
use verilog.vl_types.all;
entity ifetch is
    port(
        clock           : in     vl_logic;
        imem_address    : out    vl_logic_vector(31 downto 0);
        imem_data       : in     vl_logic_vector(127 downto 0);
        imem_read       : out    vl_logic;
        pc_address      : in     vl_logic_vector(31 downto 0);
        nxt_address     : out    vl_logic_vector(31 downto 0);
        write_pc        : out    vl_logic;
        out_op1         : out    vl_logic_vector(31 downto 0);
        out_src11       : out    vl_logic_vector(31 downto 0);
        out_src12       : out    vl_logic_vector(31 downto 0);
        out_dst1        : out    vl_logic_vector(4 downto 0);
        out_imm1        : out    vl_logic_vector(31 downto 0);
        out_srcn11      : out    vl_logic_vector(4 downto 0);
        out_srcn12      : out    vl_logic_vector(4 downto 0);
        in_src11        : in     vl_logic_vector(31 downto 0);
        in_src12        : in     vl_logic_vector(31 downto 0);
        read_src11      : out    vl_logic;
        read_src12      : out    vl_logic;
        out_op2         : out    vl_logic_vector(31 downto 0);
        out_src21       : out    vl_logic_vector(31 downto 0);
        out_src22       : out    vl_logic_vector(31 downto 0);
        out_dst2        : out    vl_logic_vector(4 downto 0);
        out_imm2        : out    vl_logic_vector(31 downto 0);
        out_srcn21      : out    vl_logic_vector(4 downto 0);
        out_srcn22      : out    vl_logic_vector(4 downto 0);
        in_src21        : in     vl_logic_vector(31 downto 0);
        in_src22        : in     vl_logic_vector(31 downto 0);
        read_src21      : out    vl_logic;
        read_src22      : out    vl_logic;
        out_op3         : out    vl_logic_vector(31 downto 0);
        out_src31       : out    vl_logic_vector(31 downto 0);
        out_src32       : out    vl_logic_vector(31 downto 0);
        out_dst3        : out    vl_logic_vector(4 downto 0);
        out_imm3        : out    vl_logic_vector(31 downto 0);
        out_srcn31      : out    vl_logic_vector(4 downto 0);
        out_srcn32      : out    vl_logic_vector(4 downto 0);
        in_src31        : in     vl_logic_vector(31 downto 0);
        in_src32        : in     vl_logic_vector(31 downto 0);
        read_src31      : out    vl_logic;
        read_src32      : out    vl_logic;
        out_op4         : out    vl_logic_vector(31 downto 0);
        out_src41       : out    vl_logic_vector(31 downto 0);
        out_src42       : out    vl_logic_vector(31 downto 0);
        out_dst4        : out    vl_logic_vector(4 downto 0);
        out_imm4        : out    vl_logic_vector(31 downto 0);
        out_srcn41      : out    vl_logic_vector(4 downto 0);
        out_srcn42      : out    vl_logic_vector(4 downto 0);
        in_src41        : in     vl_logic_vector(31 downto 0);
        in_src42        : in     vl_logic_vector(31 downto 0);
        read_src41      : out    vl_logic;
        read_src42      : out    vl_logic;
        rg_check_ok     : in     vl_logic;
        rg_check_num    : out    vl_logic_vector(4 downto 0);
        rg_check        : out    vl_logic;
        rs_op           : out    vl_logic_vector(31 downto 0);
        rs_address      : out    vl_logic_vector(31 downto 0);
        rs_reg          : out    vl_logic_vector(4 downto 0);
        rs_reg2         : out    vl_logic_vector(4 downto 0);
        rs_write        : out    vl_logic;
        rs_free         : in     vl_logic;
        rs_ex_ok        : in     vl_logic;
        in_databus      : in     vl_logic_vector(63 downto 0);
        in_databus2     : in     vl_logic_vector(63 downto 0)
    );
end ifetch;
