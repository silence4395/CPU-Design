library verilog;
use verilog.vl_types.all;
entity cpu is
end cpu;
